// $Id: $
// file_name    : NTSC_ENC.v
// descript     : for 4fsc 
//
//
//180426r       :mod for new coding rule
// 2013-02-23W6 : rename NTSC_ENC from color_enc
//                 append EE , and change more 
// 2009-07-27W1 : coding rure update
// 2004-05      : 1st.
module NTSC_ENC
(
      input             CK_i      ;
    , input tri1        XARST_i 
    , input             XR      ;
    , input             CK_EE_i      ;
    , input [ 7:0] tri0 YYs_i    
    , input [ 7:0] tri0 UUs_i    //2's  */
    , input [ 7:0] tri0 VVs_i    //2's  */
    , input        tri0 BURST_o   ; //1:BURST */
    , input        trt0 BLANK_o   ; //1:BLANK */
    , input        tri1 SYNC_o    ; //0:SYNC */
    , output[ 9:0]  VIDEOs_o ;
) ;
    reg     [ 2:0]  VIDEOs   ;
    wire    [ 2:0]  VIDEOs_a ;

    //      UU,VV is 2's s2
    reg     [ 2 :0]   YYs_D , UUs_D, VVs_D ;
    always@(posedge CK_i or negedge XARST_i) 
        if( ~ XARST_i)
        begin
            YYs_D <= 8'd0 ;
            UUs_D <= 8'd0 ;
            VVs_D <= 8'd0 ;
        end else if( CK_EE_i)
        begin
            YYs_D <= YYs_i;
            UUs_D <= UUs_i ;
            VVs_D <= VVs_i ;
        end 

    wire    [ 2 :0]  UUs_y    ;
    assign  UUs_y = ( BURST ) ? -3'd1 : (-3'd4 == UUs_d) ? -3'd3 : UUs_d ;
    wire    [ 2 :0]  VVs_y   ;
    assign  VVs_y = ( BURST ) ? 3'd0 : (-3'd4 == VVs_d) ? -3'd3 : VVs_d ;
    wire    [ 2:0]  chroma   ;
    assign  chroma = 
        (BLANK & ~ BURST) 
        ? 
            3'd0
        : (2'd0 == PHs) 
        ?
            UUs_y
        : (2'd1 == PHs) 
        ?
            VVs_y
        : (2'd2 == PHs) 
        ?
            -UUs_y
        : (2'd3 == PHs) 
        ?
            -VVs_y
        :
            3'd0
    ;
    wire    [ 2 :0]  YYs_y      ;
    assign YYs_y =
        ( ~ SYNC ) 
        ?
            3'd0
        : (BLANK | BURST) 
        ?
            3'd2
        : (YYs_d[2 :0] <= 3'd1) 
        ?
            3'd2
        :
            YYs_d[ 2 :0]
    ;

    wire    [ 4 :0]  VIDEO_aa    ;
    assign VIDEO_aa =  YYs_y + {{2{chroma[2]}} , chroma} ;
    assign VIDEO_a =
        ( ~ VIDEO_aa[ 4 ] &  VIDEO_aa[ 3 ]) 
        ?   
            3'b111
        : ( VIDEO_aa[ 4 ] ) 
        ?
            3'b000
        :
            VIDEO_aa[ 2 :0]
    ;

    always@(posedge CK_i or negedge XARST_i)
        if( ~ XARST_i )
            VIDEOs <= 10'd0 ;
        else if( CK_EE_i )
            VIDEO <= ( ~ XR) ? 3'd0 : VIDEO_a ;
    
    reg     [ 1:0]  PHs      ;  // 4fsc auto run , dont extra reset.
    always@(posedge CK_i or negedge XARST_i)
        if( ~ XARST_i)
            PHs <= 2'b0 ;
        else if( CK_EE_i )
            PHs[1:0] <= ( ~ XR) ? 2'd0 : {2{1'b1}} & (PHs + 2'd1) ;
endmodule
// NTSC_ENC.v
